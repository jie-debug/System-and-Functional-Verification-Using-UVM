class packet;
   
   //Add your code here...

endclass
