interface router_interface(input bit clk);

  //Inputs to RTL

  //Outputs from RTL

  //NOTE: The widths are 4 bits since the RTL, dut.sv, is
  //      parameterized to 4 inputs ports and 4 output ports
  //      by default. We will parameterize the interface later

  //MODPORT to indicate directions
  
endinterface
