interface switch_interface(input clk);
   //Add your code here...
endinterface
