class packet_sequence extends ...

   // Your code here

endclass
