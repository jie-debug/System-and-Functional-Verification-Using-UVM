class packet extends ...

   // Your code here

endclass

