`include "user_sequence.sv"
`include "env.sv"

class test_base extends uvm_test;

   //blah blah blah

endclass
