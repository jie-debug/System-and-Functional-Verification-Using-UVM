`include "packet.sv"

class user_sequence extends uvm_sequence #(packet);
   `uvm_object_utils(user_sequence)

endclass
