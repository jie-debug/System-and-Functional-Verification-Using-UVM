`ifndef	ENV__SV
`define	ENV__SV

`include "input_agent.sv"


class env extends uvm_env;
   `uvm_component_utils(env)

   ...
   
endclass

`endif //ENV__SV

